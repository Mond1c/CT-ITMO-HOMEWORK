package utility;
    parameter CACHE_LINE_SIZE   = 128;
    parameter CACHE_TAG_SIZE    = 8;
    parameter CACHE_SET_SIZE    = 6;
    parameter CACHE_OFFSET_SIZE = 7;



endpackage
