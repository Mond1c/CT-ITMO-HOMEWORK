module data_bus();
    parameter DATA1_BUS_SIZE = 16;
    parameter DATA2_BUS_SIZE = 16;
endmodule

module addr_bus();
    parameter ADDR1_BUS_SIZE = 14;
    parameter ADDR2_BUS_SIZE = 14;
endmodule

module ctr_bus();
    parameter CTR1_BUS_SIZE = 16;
    parameter CTR2_BUS_SIZE = 16;
endmodule;