module test;
    initial begin
        $display("Hello, world!");
    end    
endmodule